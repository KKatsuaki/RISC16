src/risc16ba.sv