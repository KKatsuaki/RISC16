geek_731@my-ubuntu.214852:1610981575