library verilog;
use verilog.vl_types.all;
entity risc16_sv_unit is
end risc16_sv_unit;
