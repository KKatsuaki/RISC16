library verilog;
use verilog.vl_types.all;
entity sim_risc16 is
end sim_risc16;
