library verilog;
use verilog.vl_types.all;
entity sim_risc16f is
end sim_risc16f;
