geek_731@MBP-KK.17402